library ieee;
use ieee.std_logic_1164.all;

entity pos_ctrl is
  port (
    -- System Clock and Reset
    rst       : in  std_logic;                    -- Reset
    rst_div   : in  std_logic;                    -- Reset
    mclk      : in  std_logic;                    -- Clock
    mclk_div  : in  std_logic;                    -- Clock to p_reg
    sync_rst  : in  std_logic;                    -- Synchronous reset
    sp        : in  std_logic_vector(7 downto 0); -- Setpoint (wanted position)
    a         : in  std_logic;                    -- From position sensor
    b         : in  std_logic;                    -- From position sensor  
    force_cw  : in  std_logic;                    -- Force motor clock wise motion
    force_ccw : in  std_logic;                    -- Force motor counter clock wise motion
    pos       : out std_logic_vector(7 downto 0); -- Measured Position
    motor_cw  : out std_logic;                    -- Motor clock wise motion
    motor_ccw : out std_logic                     -- Motor counter clock wise motion
    );      
end pos_ctrl;
